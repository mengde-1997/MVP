module top_count_32(
    input s_a0,s_a1,s_a2,s_a3,s_a4,s_a5,s_a6,s_a7,s_a8,s_a9,s_a10,s_a11,s_a12,s_a13,s_a14,s_a15,
    input s_a16,s_a17,s_a18,s_a19,s_a20,s_a21,s_a22,s_a23,s_a24,s_a25,s_a26,s_a27,s_a28,s_a29,s_a30,s_a31,
    input a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,
    input a16,a17,a18,a19,a20,a21,a22,a23,a24,a25,a26,a27,a28,a29,a30,a31,
    input [3:0]w0,w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13,w14,w15,
    input [3:0]w16,w17,w18,w19,w20,w21,w22,w23,w24,w25,w26,w27,w28,w29,w30,w31,
    output signed [15:0]h_sum
    );

    wire [6:0]h_plus_32_2,h_minus_32_2,h_plus_32_1,h_minus_32_1,h_plus_32_0,h_minus_32_0;

    assign h_sum =((h_plus_32_2-h_minus_32_2)<<2)+((h_plus_32_1-h_minus_32_1)<<1)+(h_plus_32_0-h_minus_32_0);

    count_32 count_32_2(
.t0(s_a0),.s0(w0[3]),.a0(a0),.w0(w0[2]),
.t1(s_a1),.s1(w1[3]),.a1(a1),.w1(w1[2]),
.t2(s_a2),.s2(w2[3]),.a2(a2),.w2(w2[2]),
.t3(s_a3),.s3(w3[3]),.a3(a3),.w3(w3[2]),
.t4(s_a4),.s4(w4[3]),.a4(a4),.w4(w4[2]),
.t5(s_a5),.s5(w5[3]),.a5(a5),.w5(w5[2]),
.t6(s_a6),.s6(w6[3]),.a6(a6),.w6(w6[2]),
.t7(s_a7),.s7(w7[3]),.a7(a7),.w7(w7[2]),
.t8(s_a8),.s8(w8[3]),.a8(a8),.w8(w8[2]),
.t9(s_a9),.s9(w9[3]),.a9(a9),.w9(w9[2]),
.t10(s_a10),.s10(w10[3]),.a10(a10),.w10(w10[2]),
.t11(s_a11),.s11(w11[3]),.a11(a11),.w11(w11[2]),
.t12(s_a12),.s12(w12[3]),.a12(a12),.w12(w12[2]),
.t13(s_a13),.s13(w13[3]),.a13(a13),.w13(w13[2]),
.t14(s_a14),.s14(w14[3]),.a14(a14),.w14(w14[2]),
.t15(s_a15),.s15(w15[3]),.a15(a15),.w15(w15[2]),
.t16(s_a16),.s16(w16[3]),.a16(a16),.w16(w16[2]),
.t17(s_a17),.s17(w17[3]),.a17(a17),.w17(w17[2]),
.t18(s_a18),.s18(w18[3]),.a18(a18),.w18(w18[2]),
.t19(s_a19),.s19(w19[3]),.a19(a19),.w19(w19[2]),
.t20(s_a20),.s20(w20[3]),.a20(a20),.w20(w20[2]),
.t21(s_a21),.s21(w21[3]),.a21(a21),.w21(w21[2]),
.t22(s_a22),.s22(w22[3]),.a22(a22),.w22(w22[2]),
.t23(s_a23),.s23(w23[3]),.a23(a23),.w23(w23[2]),
.t24(s_a24),.s24(w24[3]),.a24(a24),.w24(w24[2]),
.t25(s_a25),.s25(w25[3]),.a25(a25),.w25(w25[2]),
.t26(s_a26),.s26(w26[3]),.a26(a26),.w26(w26[2]),
.t27(s_a27),.s27(w27[3]),.a27(a27),.w27(w27[2]),
.t28(s_a28),.s28(w28[3]),.a28(a28),.w28(w28[2]),
.t29(s_a29),.s29(w29[3]),.a29(a29),.w29(w29[2]),
.t30(s_a30),.s30(w30[3]),.a30(a30),.w30(w30[2]),
.t31(s_a31),.s31(w31[3]),.a31(a31),.w31(w31[2]),
.h_plus_32(h_plus_32_2),.h_minus_32(h_minus_32_2)
    );

    count_32 count_32_1(
.t0(s_a0),.s0(w0[3]),.a0(a0),.w0(w0[1]),
.t1(s_a1),.s1(w1[3]),.a1(a1),.w1(w1[1]),
.t2(s_a2),.s2(w2[3]),.a2(a2),.w2(w2[1]),
.t3(s_a3),.s3(w3[3]),.a3(a3),.w3(w3[1]),
.t4(s_a4),.s4(w4[3]),.a4(a4),.w4(w4[1]),
.t5(s_a5),.s5(w5[3]),.a5(a5),.w5(w5[1]),
.t6(s_a6),.s6(w6[3]),.a6(a6),.w6(w6[1]),
.t7(s_a7),.s7(w7[3]),.a7(a7),.w7(w7[1]),
.t8(s_a8),.s8(w8[3]),.a8(a8),.w8(w8[1]),
.t9(s_a9),.s9(w9[3]),.a9(a9),.w9(w9[1]),
.t10(s_a10),.s10(w10[3]),.a10(a10),.w10(w10[1]),
.t11(s_a11),.s11(w11[3]),.a11(a11),.w11(w11[1]),
.t12(s_a12),.s12(w12[3]),.a12(a12),.w12(w12[1]),
.t13(s_a13),.s13(w13[3]),.a13(a13),.w13(w13[1]),
.t14(s_a14),.s14(w14[3]),.a14(a14),.w14(w14[1]),
.t15(s_a15),.s15(w15[3]),.a15(a15),.w15(w15[1]),
.t16(s_a16),.s16(w16[3]),.a16(a16),.w16(w16[1]),
.t17(s_a17),.s17(w17[3]),.a17(a17),.w17(w17[1]),
.t18(s_a18),.s18(w18[3]),.a18(a18),.w18(w18[1]),
.t19(s_a19),.s19(w19[3]),.a19(a19),.w19(w19[1]),
.t20(s_a20),.s20(w20[3]),.a20(a20),.w20(w20[1]),
.t21(s_a21),.s21(w21[3]),.a21(a21),.w21(w21[1]),
.t22(s_a22),.s22(w22[3]),.a22(a22),.w22(w22[1]),
.t23(s_a23),.s23(w23[3]),.a23(a23),.w23(w23[1]),
.t24(s_a24),.s24(w24[3]),.a24(a24),.w24(w24[1]),
.t25(s_a25),.s25(w25[3]),.a25(a25),.w25(w25[1]),
.t26(s_a26),.s26(w26[3]),.a26(a26),.w26(w26[1]),
.t27(s_a27),.s27(w27[3]),.a27(a27),.w27(w27[1]),
.t28(s_a28),.s28(w28[3]),.a28(a28),.w28(w28[1]),
.t29(s_a29),.s29(w29[3]),.a29(a29),.w29(w29[1]),
.t30(s_a30),.s30(w30[3]),.a30(a30),.w30(w30[1]),
.t31(s_a31),.s31(w31[3]),.a31(a31),.w31(w31[1]),
.h_plus_32(h_plus_32_1),.h_minus_32(h_minus_32_1)
    );

    count_32 count_32_0(
.t0(s_a0),.s0(w0[3]),.a0(a0),.w0(w0[0]),
.t1(s_a1),.s1(w1[3]),.a1(a1),.w1(w1[0]),
.t2(s_a2),.s2(w2[3]),.a2(a2),.w2(w2[0]),
.t3(s_a3),.s3(w3[3]),.a3(a3),.w3(w3[0]),
.t4(s_a4),.s4(w4[3]),.a4(a4),.w4(w4[0]),
.t5(s_a5),.s5(w5[3]),.a5(a5),.w5(w5[0]),
.t6(s_a6),.s6(w6[3]),.a6(a6),.w6(w6[0]),
.t7(s_a7),.s7(w7[3]),.a7(a7),.w7(w7[0]),
.t8(s_a8),.s8(w8[3]),.a8(a8),.w8(w8[0]),
.t9(s_a9),.s9(w9[3]),.a9(a9),.w9(w9[0]),
.t10(s_a10),.s10(w10[3]),.a10(a10),.w10(w10[0]),
.t11(s_a11),.s11(w11[3]),.a11(a11),.w11(w11[0]),
.t12(s_a12),.s12(w12[3]),.a12(a12),.w12(w12[0]),
.t13(s_a13),.s13(w13[3]),.a13(a13),.w13(w13[0]),
.t14(s_a14),.s14(w14[3]),.a14(a14),.w14(w14[0]),
.t15(s_a15),.s15(w15[3]),.a15(a15),.w15(w15[0]),
.t16(s_a16),.s16(w16[3]),.a16(a16),.w16(w16[0]),
.t17(s_a17),.s17(w17[3]),.a17(a17),.w17(w17[0]),
.t18(s_a18),.s18(w18[3]),.a18(a18),.w18(w18[0]),
.t19(s_a19),.s19(w19[3]),.a19(a19),.w19(w19[0]),
.t20(s_a20),.s20(w20[3]),.a20(a20),.w20(w20[0]),
.t21(s_a21),.s21(w21[3]),.a21(a21),.w21(w21[0]),
.t22(s_a22),.s22(w22[3]),.a22(a22),.w22(w22[0]),
.t23(s_a23),.s23(w23[3]),.a23(a23),.w23(w23[0]),
.t24(s_a24),.s24(w24[3]),.a24(a24),.w24(w24[0]),
.t25(s_a25),.s25(w25[3]),.a25(a25),.w25(w25[0]),
.t26(s_a26),.s26(w26[3]),.a26(a26),.w26(w26[0]),
.t27(s_a27),.s27(w27[3]),.a27(a27),.w27(w27[0]),
.t28(s_a28),.s28(w28[3]),.a28(a28),.w28(w28[0]),
.t29(s_a29),.s29(w29[3]),.a29(a29),.w29(w29[0]),
.t30(s_a30),.s30(w30[3]),.a30(a30),.w30(w30[0]),
.t31(s_a31),.s31(w31[3]),.a31(a31),.w31(w31[0]),
.h_plus_32(h_plus_32_0),.h_minus_32(h_minus_32_0)
    );

endmodule
